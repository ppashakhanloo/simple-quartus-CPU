// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 9.0 Build 132 02/25/2009 SJ Web Edition
// Created on Sun Jun 15 07:46:50 2014

// synthesis message_off 10175

`timescale 1ns/1ns

module CU (
    reset,clock,OP_4,OP_3,OP_2,OP_1,OP_0,
    COUNT_ENABLE,SEL_LOAD_PC_1,SEL_LOAD_PC_0,IR_ENABLE,SEL_AW_RF,SEL_DW_RF_1,SEL_DW_RF_0,WE_RF,SEL_IMM,SEL_INP1,SEL_INP2,SEL_ALU_3,SEL_ALU_2,SEL_ALU_1,SEL_ALU_0,WE_RAM,SEL_AR_RAM,SEL_AR2_RF);

    input reset;
    input clock;
    input OP_4;
    input OP_3;
    input OP_2;
    input OP_1;
    input OP_0;
    tri0 reset;
    tri0 OP_4;
    tri0 OP_3;
    tri0 OP_2;
    tri0 OP_1;
    tri0 OP_0;
    output COUNT_ENABLE;
    output SEL_LOAD_PC_1;
    output SEL_LOAD_PC_0;
    output IR_ENABLE;
    output SEL_AW_RF;
    output SEL_DW_RF_1;
    output SEL_DW_RF_0;
    output WE_RF;
    output SEL_IMM;
    output SEL_INP1;
    output SEL_INP2;
    output SEL_ALU_3;
    output SEL_ALU_2;
    output SEL_ALU_1;
    output SEL_ALU_0;
    output WE_RAM;
    output SEL_AR_RAM;
    output SEL_AR2_RF;
    reg COUNT_ENABLE;
    reg SEL_LOAD_PC_1;
    reg SEL_LOAD_PC_0;
    reg IR_ENABLE;
    reg SEL_AW_RF;
    reg SEL_DW_RF_1;
    reg SEL_DW_RF_0;
    reg WE_RF;
    reg SEL_IMM;
    reg SEL_INP1;
    reg SEL_INP2;
    reg SEL_ALU_3;
    reg SEL_ALU_2;
    reg SEL_ALU_1;
    reg SEL_ALU_0;
    reg WE_RAM;
    reg SEL_AR_RAM;
    reg SEL_AR2_RF;
    reg [34:0] fstate;
    reg [34:0] reg_fstate;
    parameter FETCH=0,ADD=1,SUB=2,MUL=3,DIV=4,MOD_M=5,MAX=6,MIN=7,NOT_M=8,NAND_M=9,NOR_M=10,XNOR_M=11,SHL=12,SHRA=13,ROL_M=14,ROR_M=15,LDI=16,ADDI=17,SUBI=18,MULI=19,DIVI=20,NANDI=21,NORI=22,XNORI=23,MOV=24,SWP_0=25,SWP_1=26,SWP_2=27,LD=28,STR=29,JMP=30,BEQ=31,BLT=32,HLT=33,SHRL=34;

    always @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= FETCH;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or OP_4 or OP_3 or OP_2 or OP_1 or OP_0)
    begin
        COUNT_ENABLE <= 1'b0;
        SEL_LOAD_PC_1 <= 1'b0;
        SEL_LOAD_PC_0 <= 1'b0;
        IR_ENABLE <= 1'b0;
        SEL_AW_RF <= 1'b0;
        SEL_DW_RF_1 <= 1'b0;
        SEL_DW_RF_0 <= 1'b0;
        WE_RF <= 1'b0;
        SEL_IMM <= 1'b0;
        SEL_INP1 <= 1'b0;
        SEL_INP2 <= 1'b0;
        SEL_ALU_3 <= 1'b0;
        SEL_ALU_2 <= 1'b0;
        SEL_ALU_1 <= 1'b0;
        SEL_ALU_0 <= 1'b0;
        WE_RAM <= 1'b0;
        SEL_AR_RAM <= 1'b0;
        SEL_AR2_RF <= 1'b0;
        case (fstate)
            FETCH: begin
                if ((~(OP_4) & (~(OP_3) & (~(OP_2) & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= ADD;
                else if ((~(OP_4) & (~(OP_3) & (~(OP_2) & (~(OP_1) & OP_0)))))
                    reg_fstate <= SUB;
                else if ((~(OP_4) & (~(OP_3) & (~(OP_2) & (OP_1 & ~(OP_0))))))
                    reg_fstate <= MUL;
                else if ((~(OP_4) & (~(OP_3) & (~(OP_2) & (OP_1 & OP_0)))))
                    reg_fstate <= DIV;
                else if ((~(OP_4) & (~(OP_3) & (OP_2 & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= MOD_M;
                else if ((~(OP_4) & (~(OP_3) & (OP_2 & (~(OP_1) & OP_0)))))
                    reg_fstate <= MAX;
                else if ((~(OP_4) & (~(OP_3) & (OP_2 & (OP_1 & ~(OP_0))))))
                    reg_fstate <= MIN;
                else if ((~(OP_4) & (~(OP_3) & (OP_2 & (OP_1 & OP_0)))))
                    reg_fstate <= NOT_M;
                else if ((~(OP_4) & (OP_3 & (~(OP_2) & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= NAND_M;
                else if ((~(OP_4) & (OP_3 & (~(OP_2) & (~(OP_1) & OP_0)))))
                    reg_fstate <= NOR_M;
                else if ((~(OP_4) & (OP_3 & (~(OP_2) & (OP_1 & ~(OP_0))))))
                    reg_fstate <= XNOR_M;
                else if ((~(OP_4) & (OP_3 & (~(OP_2) & (OP_1 & OP_0)))))
                    reg_fstate <= SHL;
                else if ((~(OP_4) & (OP_3 & (OP_2 & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= SHRA;
                else if ((~(OP_4) & (OP_3 & (OP_2 & (~(OP_1) & OP_0)))))
                    reg_fstate <= SHRL;
                else if ((~(OP_4) & (OP_3 & (OP_2 & (OP_1 & ~(OP_0))))))
                    reg_fstate <= ROL_M;
                else if ((~(OP_4) & (OP_3 & (OP_2 & (OP_1 & OP_0)))))
                    reg_fstate <= ROR_M;
                else if ((OP_4 & (~(OP_3) & (~(OP_2) & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= LDI;
                else if ((OP_4 & (~(OP_3) & (~(OP_2) & (~(OP_1) & OP_0)))))
                    reg_fstate <= ADDI;
                else if ((OP_4 & (~(OP_3) & (~(OP_2) & (OP_1 & ~(OP_0))))))
                    reg_fstate <= SUBI;
                else if ((OP_4 & (~(OP_3) & (~(OP_2) & (OP_1 & OP_0)))))
                    reg_fstate <= MULI;
                else if ((OP_4 & (~(OP_3) & (OP_2 & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= DIVI;
                else if ((OP_4 & (~(OP_3) & (OP_2 & (~(OP_1) & OP_0)))))
                    reg_fstate <= NANDI;
                else if ((OP_4 & (~(OP_3) & (OP_2 & (OP_1 & ~(OP_0))))))
                    reg_fstate <= NORI;
                else if ((OP_4 & (~(OP_3) & (OP_2 & (OP_1 & OP_0)))))
                    reg_fstate <= XNORI;
                else if ((OP_4 & (OP_3 & (~(OP_2) & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= MOV;
                else if ((OP_4 & (OP_3 & (~(OP_2) & (~(OP_1) & OP_0)))))
                    reg_fstate <= SWP_0;
                else if ((OP_4 & (OP_3 & (~(OP_2) & (OP_1 & ~(OP_0))))))
                    reg_fstate <= LD;
                else if ((OP_4 & (OP_3 & (~(OP_2) & (OP_1 & OP_0)))))
                    reg_fstate <= STR;
                else if ((OP_4 & (OP_3 & (OP_2 & (~(OP_1) & ~(OP_0))))))
                    reg_fstate <= JMP;
                else if ((OP_4 & (OP_3 & (OP_2 & (~(OP_1) & OP_0)))))
                    reg_fstate <= BEQ;
                else if ((OP_4 & (OP_3 & (OP_2 & (OP_1 & ~(OP_0))))))
                    reg_fstate <= BLT;
                else if ((OP_4 & (OP_3 & (OP_2 & (OP_1 & OP_0)))))
                    reg_fstate <= HLT;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b0;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b1;

                WE_RF <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR_RAM <= 1'b0;
            end
            ADD: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            SUB: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            MUL: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            DIV: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            MOD_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            MAX: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            MIN: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            NOT_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            NAND_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            NOR_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            XNOR_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b1;
            end
            SHL: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            SHRA: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            ROL_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            ROR_M: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            LDI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b0;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            ADDI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            SUBI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            MULI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            DIVI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            NANDI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            NORI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            XNORI: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b1;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            MOV: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_IMM <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b1;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;
            end
            SWP_0: begin
                reg_fstate <= SWP_1;

                COUNT_ENABLE <= 1'b0;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                WE_RF <= 1'b0;

                WE_RAM <= 1'b0;
            end
            SWP_1: begin
                reg_fstate <= SWP_2;

                COUNT_ENABLE <= 1'b0;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b1;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b0;

                SEL_INP2 <= 1'b0;

                SEL_ALU_3 <= 1'b0;

                SEL_ALU_2 <= 1'b0;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b0;
            end
            SWP_2: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b1;

                SEL_DW_RF_0 <= 1'b0;

                WE_RF <= 1'b1;

                WE_RAM <= 1'b0;
            end
            LD: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b0;

                WE_RF <= 1'b1;

                WE_RAM <= 1'b0;

                SEL_AR_RAM <= 1'b1;
            end
            STR: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                WE_RF <= 1'b0;

                SEL_INP2 <= 1'b0;

                WE_RAM <= 1'b1;

                SEL_AR_RAM <= 1'b1;

                SEL_AR2_RF <= 1'b0;
            end
            JMP: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b0;

                SEL_LOAD_PC_0 <= 1'b0;

                IR_ENABLE <= 1'b0;

                WE_RF <= 1'b0;

                WE_RAM <= 1'b0;
            end
            BEQ: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b0;

                IR_ENABLE <= 1'b0;

                WE_RF <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b0;
            end
            BLT: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b0;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                WE_RF <= 1'b0;

                SEL_INP1 <= 1'b1;

                SEL_INP2 <= 1'b0;

                WE_RAM <= 1'b0;

                SEL_AR2_RF <= 1'b0;
            end
            HLT: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b0;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                WE_RF <= 1'b0;

                WE_RAM <= 1'b0;
            end
            SHRL: begin
                reg_fstate <= FETCH;

                COUNT_ENABLE <= 1'b1;

                SEL_LOAD_PC_1 <= 1'b1;

                SEL_LOAD_PC_0 <= 1'b1;

                IR_ENABLE <= 1'b0;

                SEL_AW_RF <= 1'b0;

                SEL_DW_RF_1 <= 1'b0;

                SEL_DW_RF_0 <= 1'b1;

                WE_RF <= 1'b1;

                SEL_INP1 <= 1'b1;

                SEL_ALU_3 <= 1'b1;

                SEL_ALU_2 <= 1'b1;

                SEL_ALU_1 <= 1'b0;

                SEL_ALU_0 <= 1'b1;

                WE_RAM <= 1'b0;
            end
            default: begin
                COUNT_ENABLE <= 1'bx;
                SEL_LOAD_PC_1 <= 1'bx;
                SEL_LOAD_PC_0 <= 1'bx;
                IR_ENABLE <= 1'bx;
                SEL_AW_RF <= 1'bx;
                SEL_DW_RF_1 <= 1'bx;
                SEL_DW_RF_0 <= 1'bx;
                WE_RF <= 1'bx;
                SEL_IMM <= 1'bx;
                SEL_INP1 <= 1'bx;
                SEL_INP2 <= 1'bx;
                SEL_ALU_3 <= 1'bx;
                SEL_ALU_2 <= 1'bx;
                SEL_ALU_1 <= 1'bx;
                SEL_ALU_0 <= 1'bx;
                WE_RAM <= 1'bx;
                SEL_AR_RAM <= 1'bx;
                SEL_AR2_RF <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // CU

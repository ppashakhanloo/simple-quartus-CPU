module MEMORY (DATA_OUT, DATA_IN, ADDRESS_READ, ADDRESS_WRITE, CLK, RESET, WRITE_ENABLE);
  
  output [31 : 0] DATA_OUT;
  input [31 : 0] DATA_IN;
  input [7 : 0] ADDRESS_READ, ADDRESS_WRITE;
  input CLK, RESET, WRITE_ENABLE;
  
  reg [31 : 0] Memory [0 : 255];
  
  assign DATA_OUT = Memory [ADDRESS_READ];
  
  always @(posedge CLK or posedge RESET)
    if (RESET)  begin
      //Your code goes here.
      Memory [000] = 32'b10000000010000000000000000000010;	// $1 <- 1	
      Memory [001] = 32'b10000000100000000000000000000100;	// $2 <- 2
      Memory [002] = 32'b00010000000000100010000000000000;	// $0 <- $1 * $2
      Memory [003] = 32'b10000000110000000000000000000110;	// $3 <- 3
      Memory [004] = 32'b10000000110000000000000000010110;	// $3 <- 11	
      Memory [005] = 32'b11010000000000100000000000000000;	// 	
      Memory [006] = 32'b11011000100001100000000000000000;	//	
      Memory [007] = 32'b11010000010001100000000000000000;	// 
      Memory [008] = 32'b11111000010000100000000000000100;	// 	
      Memory [009] = 32'b11111000000000000000000000000000;	// halt
      Memory [010] = 32'b00000000000000000000000000000000;		
      Memory [011] = 32'b01010101010101010101010101010101;		
      Memory [012] = 32'b00000000000000000000000000000000;			
      Memory [013] = 32'b00000000000000000000000000000000;			
      Memory [014] = 32'b00000000000000000000000000000000;			
      Memory [015] = 32'b00000000000000000000000000000000;			
      Memory [016] = 32'b00000000000000000000000000000000;			
      Memory [017] = 32'b00000000000000000000000000000000;		
      Memory [018] = 32'b00000000000000000000000000000000;		
      Memory [019] = 32'b00000000000000000000000000000000;		
      Memory [020] = 32'b00000000000000000000000000000000;		
      Memory [021] = 32'b00000000000000000000000000000000;		
      Memory [022] = 32'b00000000000000000000000000000000;		
      Memory [023] = 32'b00000000000000000000000000000000;
      Memory [024] = 32'b00000000000000000000000000000000;
      Memory [025] = 32'b00000000000000000000000000000000;
      Memory [026] = 32'b00000000000000000000000000000000;
      Memory [027] = 32'b00000000000000000000000000000000;
      Memory [028] = 32'b00000000000000000000000000000000;
      Memory [029] = 32'b00000000000000000000000000000000;
      Memory [030] = 32'b00000000000000000000000000000000;
      Memory [031] = 32'b00000000000000000000000000000000;			
      Memory [032] = 32'b00000000000000000000000000000000;			
      Memory [033] = 32'b00000000000000000000000000000000;
      Memory [034] = 32'b00000000000000000000000000000000;
      Memory [035] = 32'b00000000000000000000000000000000;
      Memory [036] = 32'b00000000000000000000000000000000;
      Memory [037] = 32'b00000000000000000000000000000000;
      Memory [038] = 32'b00000000000000000000000000000000;
      Memory [039] = 32'b00000000000000000000000000000000;
      Memory [040] = 32'b00000000000000000000000000000000;
      Memory [041] = 32'b00000000000000000000000000000000;
      Memory [042] = 32'b00000000000000000000000000000000;
      Memory [043] = 32'b00000000000000000000000000000000;
      Memory [044] = 32'b00000000000000000000000000000000;
      Memory [045] = 32'b00000000000000000000000000000000;
      Memory [046] = 32'b00000000000000000000000000000000;
      Memory [047] = 32'b00000000000000000000000000000000;
      Memory [048] = 32'b00000000000000000000000000000000;
      Memory [049] = 32'b00000000000000000000000000000000;
      Memory [050] = 32'b00000000000000000000000000000000;
      Memory [051] = 32'b00000000000000000000000000000000;
      Memory [052] = 32'b00000000000000000000000000000000;
      Memory [053] = 32'b00000000000000000000000000000000;
      Memory [054] = 32'b00000000000000000000000000000000;
      Memory [055] = 32'b00000000000000000000000000000000;
      Memory [056] = 32'b00000000000000000000000000000000;
      Memory [057] = 32'b00000000000000000000000000000000;
      Memory [058] = 32'b00000000000000000000000000000000;
      Memory [059] = 32'b00000000000000000000000000000000;
      Memory [060] = 32'b00000000000000000000000000000000;
      Memory [061] = 32'b00000000000000000000000000000000;
      Memory [062] = 32'b00000000000000000000000000000000;
      Memory [063] = 32'b00000000000000000000000000000000;
      Memory [064] = 32'b00000000000000000000000000000000;
      Memory [065] = 32'b00000000000000000000000000000000;
      Memory [066] = 32'b00000000000000000000000000000000;
      Memory [067] = 32'b00000000000000000000000000000000;
      Memory [068] = 32'b00000000000000000000000000000000;
      Memory [069] = 32'b00000000000000000000000000000000;
      Memory [070] = 32'b00000000000000000000000000000000;
      Memory [071] = 32'b00000000000000000000000000000000;
      Memory [072] = 32'b00000000000000000000000000000000;
      Memory [073] = 32'b00000000000000000000000000000000;
      Memory [074] = 32'b00000000000000000000000000000000;
      Memory [075] = 32'b00000000000000000000000000000000;
      Memory [076] = 32'b00000000000000000000000000000000;
      Memory [077] = 32'b00000000000000000000000000000000;
      Memory [078] = 32'b00000000000000000000000000000000;
      Memory [079] = 32'b00000000000000000000000000000000;
      Memory [080] = 32'b00000000000000000000000000000000;
      Memory [081] = 32'b00000000000000000000000000000000;
      Memory [082] = 32'b00000000000000000000000000000000;
      Memory [083] = 32'b00000000000000000000000000000000;
      Memory [084] = 32'b00000000000000000000000000000000;
      Memory [085] = 32'b00000000000000000000000000000000;
      Memory [086] = 32'b00000000000000000000000000000000;
      Memory [087] = 32'b00000000000000000000000000000000;
      Memory [088] = 32'b00000000000000000000000000000000;
      Memory [089] = 32'b00000000000000000000000000000000;
      Memory [090] = 32'b00000000000000000000000000000000;
      Memory [091] = 32'b00000000000000000000000000000000;
      Memory [092] = 32'b00000000000000000000000000000000;
      Memory [093] = 32'b00000000000000000000000000000000;
      Memory [094] = 32'b00000000000000000000000000000000;
      Memory [095] = 32'b00000000000000000000000000000000;
      Memory [096] = 32'b00000000000000000000000000000000;
      Memory [097] = 32'b00000000000000000000000000000000;
      Memory [098] = 32'b00000000000000000000000000000000;
      Memory [099] = 32'b00000000000000000000000000000000;
      Memory [100] = 32'b00000000000000000000000000000000;
      Memory [101] = 32'b00000000000000000000000000000000;
      Memory [102] = 32'b00000000000000000000000000000000;
      Memory [103] = 32'b00000000000000000000000000000000;
      Memory [104] = 32'b00000000000000000000000000000000;
      Memory [105] = 32'b00000000000000000000000000000000;
      Memory [106] = 32'b00000000000000000000000000000000;
      Memory [107] = 32'b00000000000000000000000000000000;
      Memory [108] = 32'b00000000000000000000000000000000;
      Memory [109] = 32'b00000000000000000000000000000000;
      Memory [110] = 32'b00000000000000000000000000000000;
      Memory [111] = 32'b00000000000000000000000000000000;
      Memory [112] = 32'b00000000000000000000000000000000;
      Memory [113] = 32'b00000000000000000000000000000000;
      Memory [114] = 32'b00000000000000000000000000000000;
      Memory [115] = 32'b00000000000000000000000000000000;
      Memory [116] = 32'b00000000000000000000000000000000;
      Memory [117] = 32'b00000000000000000000000000000000;
      Memory [118] = 32'b00000000000000000000000000000000;
      Memory [119] = 32'b00000000000000000000000000000000;
      Memory [120] = 32'b00000000000000000000000000000000;
      Memory [121] = 32'b00000000000000000000000000000000;
      Memory [122] = 32'b00000000000000000000000000000000;
      Memory [123] = 32'b00000000000000000000000000000000;
      Memory [124] = 32'b00000000000000000000000000000000;
      Memory [125] = 32'b00000000000000000000000000000000;
      Memory [126] = 32'b00000000000000000000000000000000;
      Memory [127] = 32'b00000000000000000000000000000000;
      Memory [128] = 32'b00000000000000000000000000000000;
      Memory [129] = 32'b00000000000000000000000000000000;
      Memory [130] = 32'b00000000000000000000000000000000;
      Memory [131] = 32'b00000000000000000000000000000000;
      Memory [132] = 32'b00000000000000000000000000000000;
      Memory [133] = 32'b00000000000000000000000000000000;
      Memory [134] = 32'b00000000000000000000000000000000;
      Memory [135] = 32'b00000000000000000000000000000000;
      Memory [136] = 32'b00000000000000000000000000000000;
      Memory [137] = 32'b00000000000000000000000000000000;
      Memory [138] = 32'b00000000000000000000000000000000;
      Memory [139] = 32'b00000000000000000000000000000000;
      Memory [140] = 32'b00000000000000000000000000000000;
      Memory [141] = 32'b00000000000000000000000000000000;
      Memory [142] = 32'b00000000000000000000000000000000;
      Memory [143] = 32'b00000000000000000000000000000000;
      Memory [144] = 32'b00000000000000000000000000000000;
      Memory [145] = 32'b00000000000000000000000000000000;
      Memory [146] = 32'b00000000000000000000000000000000;
      Memory [147] = 32'b00000000000000000000000000000000;
      Memory [148] = 32'b00000000000000000000000000000000;
      Memory [149] = 32'b00000000000000000000000000000000;
      Memory [150] = 32'b00000000000000000000000000000000;
      Memory [151] = 32'b00000000000000000000000000000000;
      Memory [152] = 32'b00000000000000000000000000000000;
      Memory [153] = 32'b00000000000000000000000000000000;
      Memory [154] = 32'b00000000000000000000000000000000;
      Memory [155] = 32'b00000000000000000000000000000000;
      Memory [156] = 32'b00000000000000000000000000000000;
      Memory [157] = 32'b00000000000000000000000000000000;
      Memory [158] = 32'b00000000000000000000000000000000;
      Memory [159] = 32'b00000000000000000000000000000000;
      Memory [160] = 32'b00000000000000000000000000000000;
      Memory [161] = 32'b00000000000000000000000000000000;
      Memory [162] = 32'b00000000000000000000000000000000;
      Memory [163] = 32'b00000000000000000000000000000000;
      Memory [164] = 32'b00000000000000000000000000000000;
      Memory [165] = 32'b00000000000000000000000000000000;
      Memory [166] = 32'b00000000000000000000000000000000;
      Memory [167] = 32'b00000000000000000000000000000000;
      Memory [168] = 32'b00000000000000000000000000000000;
      Memory [169] = 32'b00000000000000000000000000000000;
      Memory [170] = 32'b00000000000000000000000000000000;
      Memory [171] = 32'b00000000000000000000000000000000;
      Memory [172] = 32'b00000000000000000000000000000000;
      Memory [173] = 32'b00000000000000000000000000000000;
      Memory [174] = 32'b00000000000000000000000000000000;
      Memory [175] = 32'b00000000000000000000000000000000;
      Memory [176] = 32'b00000000000000000000000000000000;
      Memory [177] = 32'b00000000000000000000000000000000;
      Memory [178] = 32'b00000000000000000000000000000000;
      Memory [179] = 32'b00000000000000000000000000000000;
      Memory [180] = 32'b00000000000000000000000000000000;
      Memory [181] = 32'b00000000000000000000000000000000;
      Memory [182] = 32'b00000000000000000000000000000000;
      Memory [183] = 32'b00000000000000000000000000000000;
      Memory [184] = 32'b00000000000000000000000000000000;
      Memory [185] = 32'b00000000000000000000000000000000;
      Memory [186] = 32'b00000000000000000000000000000000;
      Memory [187] = 32'b00000000000000000000000000000000;
      Memory [188] = 32'b00000000000000000000000000000000;
      Memory [189] = 32'b00000000000000000000000000000000;
      Memory [190] = 32'b00000000000000000000000000000000;
      Memory [191] = 32'b00000000000000000000000000000000;
      Memory [192] = 32'b00000000000000000000000000000000;
      Memory [193] = 32'b00000000000000000000000000000000;
      Memory [194] = 32'b00000000000000000000000000000000;
      Memory [195] = 32'b00000000000000000000000000000000;
      Memory [196] = 32'b00000000000000000000000000000000;
      Memory [197] = 32'b00000000000000000000000000000000;
      Memory [198] = 32'b00000000000000000000000000000000;
      Memory [199] = 32'b00000000000000000000000000000000;
      Memory [200] = 32'b00000000000000000000000000000000;
      Memory [201] = 32'b00000000000000000000000000000000;
      Memory [202] = 32'b00000000000000000000000000000000;
      Memory [203] = 32'b00000000000000000000000000000000;
      Memory [204] = 32'b00000000000000000000000000000000;
      Memory [205] = 32'b00000000000000000000000000000000;
      Memory [206] = 32'b00000000000000000000000000000000;
      Memory [207] = 32'b00000000000000000000000000000000;
      Memory [208] = 32'b00000000000000000000000000000000;
      Memory [209] = 32'b00000000000000000000000000000000;
      Memory [210] = 32'b00000000000000000000000000000000;
      Memory [211] = 32'b00000000000000000000000000000000;
      Memory [212] = 32'b00000000000000000000000000000000;
      Memory [213] = 32'b00000000000000000000000000000000;
      Memory [214] = 32'b00000000000000000000000000000000;
      Memory [215] = 32'b00000000000000000000000000000000;
      Memory [216] = 32'b00000000000000000000000000000000;
      Memory [217] = 32'b00000000000000000000000000000000;
      Memory [218] = 32'b00000000000000000000000000000000;
      Memory [219] = 32'b00000000000000000000000000000000;
      Memory [220] = 32'b00000000000000000000000000000000;
      Memory [221] = 32'b00000000000000000000000000000000;
      Memory [222] = 32'b00000000000000000000000000000000;
      Memory [223] = 32'b00000000000000000000000000000000;
      Memory [224] = 32'b00000000000000000000000000000000;
      Memory [225] = 32'b00000000000000000000000000000000;
      Memory [226] = 32'b00000000000000000000000000000000;
      Memory [227] = 32'b00000000000000000000000000000000;
      Memory [228] = 32'b00000000000000000000000000000000;
      Memory [229] = 32'b00000000000000000000000000000000;
      Memory [230] = 32'b00000000000000000000000000000000;
      Memory [231] = 32'b00000000000000000000000000000000;
      Memory [232] = 32'b00000000000000000000000000000000;
      Memory [233] = 32'b00000000000000000000000000000000;
      Memory [234] = 32'b00000000000000000000000000000000;
      Memory [235] = 32'b00000000000000000000000000000000;
      Memory [236] = 32'b00000000000000000000000000000000;
      Memory [237] = 32'b00000000000000000000000000000000;
      Memory [238] = 32'b00000000000000000000000000000000;
      Memory [239] = 32'b00000000000000000000000000000000;
      Memory [240] = 32'b00000000000000000000000000000000;
      Memory [241] = 32'b00000000000000000000000000000000;
      Memory [242] = 32'b00000000000000000000000000000000;
      Memory [243] = 32'b00000000000000000000000000000000;
      Memory [244] = 32'b00000000000000000000000000000000;
      Memory [245] = 32'b00000000000000000000000000000000;
      Memory [246] = 32'b00000000000000000000000000000000;
      Memory [247] = 32'b00000000000000000000000000000000;
      Memory [248] = 32'b00000000000000000000000000000000;
      Memory [249] = 32'b00000000000000000000000000000000;
      Memory [250] = 32'b00000000000000000000000000000000;
      Memory [251] = 32'b00000000000000000000000000000000;
      Memory [252] = 32'b00000000000000000000000000000000;
      Memory [253] = 32'b00000000000000000000000000000000;
      Memory [254] = 32'b00000000000000000000000000000000;
      Memory [255] = 32'b00000000000000000000000000000000;  
    end else  if (WRITE_ENABLE)
      Memory [ADDRESS_WRITE] = DATA_IN;
    
endmodule


-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 132 02/25/2009 SJ Web Edition
-- Created on Tue Jun 10 06:14:20 2014

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CU IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        OP_4 : IN STD_LOGIC := '0';
        OP_3 : IN STD_LOGIC := '0';
        OP_2 : IN STD_LOGIC := '0';
        OP_1 : IN STD_LOGIC := '0';
        OP_0 : IN STD_LOGIC := '0';
        COUNT_ENABLE : OUT STD_LOGIC;
        SEL_LOAD_PC_1 : OUT STD_LOGIC;
        SEL_LOAD_PC_0 : OUT STD_LOGIC;
        IR_ENABLE_SEL_AR_RAM : OUT STD_LOGIC;
        SEL_AW_RF_SEL_AR2_RF : OUT STD_LOGIC;
        SEL_DW_RF_1 : OUT STD_LOGIC;
        SEL_DW_RF_0 : OUT STD_LOGIC;
        WE_RF : OUT STD_LOGIC;
        SEL_IMM : OUT STD_LOGIC;
        SEL_INP1 : OUT STD_LOGIC;
        SEL_INP2 : OUT STD_LOGIC;
        SEL_ALU_3 : OUT STD_LOGIC;
        SEL_ALU_2 : OUT STD_LOGIC;
        SEL_ALU_1 : OUT STD_LOGIC;
        SEL_ALU_0 : OUT STD_LOGIC;
        WE_RAM : OUT STD_LOGIC
    );
END CU;

ARCHITECTURE BEHAVIOR OF CU IS
    TYPE type_fstate IS (FETCH,ADD,SUB,MUL,DIV,MOD_M,MAX,MIN,NOT_M,NAND_M,NOR_M,XNOR_M,SHL,SHRA,ROL_M,ROR_M,LDI,ADDI,SUBI,MULI,DIVI,NANDI,NORI,XNORI,MOV,SWP_0,SWP_1,SWP_2,LD,STR,JMP,BEQ,BLT,HLT,SHRL);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,OP_4,OP_3,OP_2,OP_1,OP_0)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= FETCH;
            COUNT_ENABLE <= '0';
            SEL_LOAD_PC_1 <= '0';
            SEL_LOAD_PC_0 <= '0';
            IR_ENABLE_SEL_AR_RAM <= '0';
            SEL_AW_RF_SEL_AR2_RF <= '0';
            SEL_DW_RF_1 <= '0';
            SEL_DW_RF_0 <= '0';
            WE_RF <= '0';
            SEL_IMM <= '0';
            SEL_INP1 <= '0';
            SEL_INP2 <= '0';
            SEL_ALU_3 <= '0';
            SEL_ALU_2 <= '0';
            SEL_ALU_1 <= '0';
            SEL_ALU_0 <= '0';
            WE_RAM <= '0';
        ELSE
            COUNT_ENABLE <= '0';
            SEL_LOAD_PC_1 <= '0';
            SEL_LOAD_PC_0 <= '0';
            IR_ENABLE_SEL_AR_RAM <= '0';
            SEL_AW_RF_SEL_AR2_RF <= '0';
            SEL_DW_RF_1 <= '0';
            SEL_DW_RF_0 <= '0';
            WE_RF <= '0';
            SEL_IMM <= '0';
            SEL_INP1 <= '0';
            SEL_INP2 <= '0';
            SEL_ALU_3 <= '0';
            SEL_ALU_2 <= '0';
            SEL_ALU_1 <= '0';
            SEL_ALU_0 <= '0';
            WE_RAM <= '0';
            CASE fstate IS
                WHEN FETCH =>
                    IF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= ADD;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= SUB;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= MUL;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= DIV;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= MOD_M;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= MAX;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= MIN;
                    ELSIF ((NOT((OP_4 = '1')) AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= NOT_M;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= NAND_M;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= NOR_M;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= XNOR_M;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= SHL;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= SHRA;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= SHRL;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND ((OP_2 = '1') AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= ROL_M;
                    ELSIF ((NOT((OP_4 = '1')) AND ((OP_3 = '1') AND ((OP_2 = '1') AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= ROR_M;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= LDI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= ADDI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= SUBI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= MULI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= DIVI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= NANDI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= NORI;
                    ELSIF (((OP_4 = '1') AND (NOT((OP_3 = '1')) AND ((OP_2 = '1') AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= XNORI;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= MOV;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= SWP_0;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= LD;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND (NOT((OP_2 = '1')) AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= STR;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= JMP;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND ((OP_2 = '1') AND (NOT((OP_1 = '1')) AND (OP_0 = '1')))))) THEN
                        reg_fstate <= BEQ;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND ((OP_2 = '1') AND ((OP_1 = '1') AND NOT((OP_0 = '1'))))))) THEN
                        reg_fstate <= BLT;
                    ELSIF (((OP_4 = '1') AND ((OP_3 = '1') AND ((OP_2 = '1') AND ((OP_1 = '1') AND (OP_0 = '1')))))) THEN
                        reg_fstate <= HLT;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= FETCH;
                    END IF;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '1';

                    WE_RF <= '0';

                    WE_RAM <= '0';
                WHEN ADD =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN SUB =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN MUL =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN DIV =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN MOD_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN MAX =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN MIN =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN NOT_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN NAND_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN NOR_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN XNOR_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN SHL =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN SHRA =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN ROL_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN ROR_M =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN LDI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '0';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN ADDI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN SUBI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN MULI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN DIVI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN NANDI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN NORI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN XNORI =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '1';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN MOV =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_IMM <= '1';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '1';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN SWP_0 =>
                    reg_fstate <= SWP_1;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    WE_RF <= '0';

                    WE_RAM <= '0';
                WHEN SWP_1 =>
                    reg_fstate <= SWP_2;

                    COUNT_ENABLE <= '0';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '1';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '0';

                    SEL_INP2 <= '0';

                    SEL_ALU_3 <= '0';

                    SEL_ALU_2 <= '0';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '0';

                    WE_RAM <= '0';
                WHEN SWP_2 =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '0';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '1';

                    SEL_DW_RF_0 <= '0';

                    WE_RF <= '1';

                    WE_RAM <= '0';
                WHEN LD =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '0';

                    WE_RF <= '1';

                    WE_RAM <= '0';
                WHEN STR =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    WE_RF <= '0';

                    SEL_INP2 <= '0';

                    WE_RAM <= '1';
                WHEN JMP =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '0';

                    SEL_LOAD_PC_0 <= '0';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    WE_RF <= '0';

                    WE_RAM <= '0';
                WHEN BEQ =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '0';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    WE_RF <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    WE_RAM <= '0';
                WHEN BLT =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '0';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    WE_RF <= '0';

                    SEL_INP1 <= '1';

                    SEL_INP2 <= '0';

                    WE_RAM <= '0';
                WHEN HLT =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '0';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    WE_RF <= '0';

                    WE_RAM <= '0';
                WHEN SHRL =>
                    reg_fstate <= FETCH;

                    COUNT_ENABLE <= '1';

                    SEL_LOAD_PC_1 <= '1';

                    SEL_LOAD_PC_0 <= '1';

                    IR_ENABLE_SEL_AR_RAM <= '0';

                    SEL_AW_RF_SEL_AR2_RF <= '0';

                    SEL_DW_RF_1 <= '0';

                    SEL_DW_RF_0 <= '1';

                    WE_RF <= '1';

                    SEL_INP1 <= '1';

                    SEL_ALU_3 <= '1';

                    SEL_ALU_2 <= '1';

                    SEL_ALU_1 <= '0';

                    SEL_ALU_0 <= '1';

                    WE_RAM <= '0';
                WHEN OTHERS => 
                    COUNT_ENABLE <= 'X';
                    SEL_LOAD_PC_1 <= 'X';
                    SEL_LOAD_PC_0 <= 'X';
                    IR_ENABLE_SEL_AR_RAM <= 'X';
                    SEL_AW_RF_SEL_AR2_RF <= 'X';
                    SEL_DW_RF_1 <= 'X';
                    SEL_DW_RF_0 <= 'X';
                    WE_RF <= 'X';
                    SEL_IMM <= 'X';
                    SEL_INP1 <= 'X';
                    SEL_INP2 <= 'X';
                    SEL_ALU_3 <= 'X';
                    SEL_ALU_2 <= 'X';
                    SEL_ALU_1 <= 'X';
                    SEL_ALU_0 <= 'X';
                    WE_RAM <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
